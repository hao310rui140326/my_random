module test_case();


endmodule


